library verilog;
use verilog.vl_types.all;
entity DiceTest_vlg_vec_tst is
end DiceTest_vlg_vec_tst;
